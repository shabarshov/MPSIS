module inv (
    input logic A,
    output logic D
);

assign D = ~A;

endmodule